-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.0 Build 156 04/24/2013 SJ Web Edition"
-- CREATED		"Thu Sep 17"
-- AUTHOR 		Bultot Geoffrey
-- LICENSE 		All right reserved

-- CE COMPOSANT PREND EN ENTREE UNE VALEUR ENTRE 0 ET 4095 VENANT D UN CAPTEUR sharp 0a41sk Et donne sa mesure sur 4 digits (dizaines, unités, dixièmes, centièmes)

-- fréquence de rafraichissement de la mesure en sortie : 2HZ

LIBRARY ieee;
USE ieee.std_logic_1164.all; 
use ieee.numeric_std.all;
use ieee.math_real.all;

LIBRARY work;

ENTITY rawTo4Digit IS 
	PORT
	(
		-- clock (50MHZ en entrée
		CLOCK_50MHZ : in std_logic;
		-- Valeur d'entrée sur 12 bits (ADC 12BITS)
		RAW_VALUE_IN : in std_logic_vector (11 downto 0);
		-- Digits de sortie sur 4 bits
		DigitDecade : out std_logic_vector (3 downto 0);
		DigitUnit : out std_logic_vector (3 downto 0);
		DigitTenth : out std_logic_vector (3 downto 0);
		DigitHundredth : out std_logic_vector (3 downto 0)
	);
END rawTo4Digit;


--*************************************************************************************
--**************** ARCHITECTURE Behavioral OF rawTo4Digit *****************************
--*************************************************************************************

ARCHITECTURE Behavioral OF rawTo4Digit IS 

-- signal clock divided (5Hz) to refresh digits
signal sig_refreshDigits : std_logic := '0';

-- Variables pour diviser la fréquence pour l'affichage des digits
shared variable temp : integer := 12499999;

BEGIN 
	-- process to divide clock in order to refresh digits 
	process(CLOCK_50MHZ)
		begin
			if rising_edge(CLOCK_50MHZ) then
				temp := temp + 1;
				if (temp=12500000) then -- 50MHZ/2/2hz = 12 500 000 (divise par 2 parce que rising_edge)
					-- frequence divided
					sig_refreshDigits <= not(sig_refreshDigits);
					temp:=0; 
				end if;
			end if;
		end process;


	refreshOutput : process(sig_refreshDigits)
		variable realValue : integer := 0;
		begin
			if falling_edge(sig_refreshDigits) then
					-- Conversion. see sensor datasheet for more informations
					realValue := 717144 / (to_integer(unsigned(RAW_VALUE_IN))/2);-- 13 * 4096 * 100 / (RAW*VOLTAGE(5)) 
					--4096/5V : 1064960 
					--2048/5V : 532480  
					--4096/3V3 : 1613575 CORRIG(/9*8) : 1434288
					--2048/3V3 : 806787 CORRIG(/9*8) : 717144
					
					--uncomment to have raw value to digits
					--realValue := to_integer(unsigned(RAW_VALUE_IN));
					
					DigitHundredth  <= std_logic_vector(to_unsigned(realValue mod 10, DigitHundredth'length));
					realValue := realValue/10;
					DigitTenth<= std_logic_vector(to_unsigned((realValue) mod 10, DigitTenth'length));
					realValue := realValue/10;
					DigitUnit  <= std_logic_vector(to_unsigned((realValue) mod 10, DigitUnit'length));
					realValue := realValue/10;
					DigitDecade<= std_logic_vector(to_unsigned((realValue) mod 10, DigitDecade'length));
			end if;
		end process;
END Behavioral;

